library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity camera is
  port (
    clock
  ) ;
end camera ;

architecture arch of camera is



begin



end architecture ; -- arch